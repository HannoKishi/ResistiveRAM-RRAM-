module decoder_5to32(en,din,dout);
 input en;
 input [4:0] din;
 output[31:0] dout;
 reg [31:0] dout;
 always@(din or en)
  begin
   if(!en)
    dout=0;
   else 
    case(din)
	 5'b00000: dout=32'b0000_0000_0000_0000_0000_0000_0000_0001;
	 5'b00001: dout=32'b0000_0000_0000_0000_0000_0000_0000_0010;
	 5'b00010: dout=32'b0000_0000_0000_0000_0000_0000_0000_0100;
	 5'b00011: dout=32'b0000_0000_0000_0000_0000_0000_0000_1000;
	 5'b00100: dout=32'b0000_0000_0000_0000_0000_0000_0001_0000;
	 5'b00101: dout=32'b0000_0000_0000_0000_0000_0000_0010_0000;
	 5'b00110: dout=32'b0000_0000_0000_0000_0000_0000_0100_0000;
	 5'b00111: dout=32'b0000_0000_0000_0000_0000_0000_1000_0000;
	 5'b01000: dout=32'b0000_0000_0000_0000_0000_0001_0000_0000;
	 5'b01001: dout=32'b0000_0000_0000_0000_0000_0010_0000_0000;
	 5'b01010: dout=32'b0000_0000_0000_0000_0000_0100_0000_0000;
	 5'b01011: dout=32'b0000_0000_0000_0000_0000_1000_0000_0000;
	 5'b01100: dout=32'b0000_0000_0000_0000_0001_0000_0000_0000;
	 5'b01101: dout=32'b0000_0000_0000_0000_0010_0000_0000_0000;
	 5'b01110: dout=32'b0000_0000_0000_0000_0100_0000_0000_0000;
	 5'b01111: dout=32'b0000_0000_0000_0000_1000_0000_0000_0000;
	 5'b10000: dout=32'b0000_0000_0000_0001_0000_0000_0000_0000;
	 5'b10001: dout=32'b0000_0000_0000_0010_0000_0000_0000_0000;
	 5'b10010: dout=32'b0000_0000_0000_0100_0000_0000_0000_0000;
	 5'b10011: dout=32'b0000_0000_0000_1000_0000_0000_0000_0000;
	 5'b10100: dout=32'b0000_0000_0001_0000_0000_0000_0000_0000;
	 5'b10101: dout=32'b0000_0000_0010_0000_0000_0000_0000_0000;
	 5'b10110: dout=32'b0000_0000_0100_0000_0000_0000_0000_0000;
	 5'b10111: dout=32'b0000_0000_1000_0000_0000_0000_0000_0000;
	 5'b11000: dout=32'b0000_0001_0000_0000_0000_0000_0000_0000;
	 5'b11001: dout=32'b0000_0010_0000_0000_0000_0000_0000_0000;
	 5'b11010: dout=32'b0000_0100_0000_0000_0000_0000_0000_0000;
	 5'b11011: dout=32'b0000_1000_0000_0000_0000_0000_0000_0000;
	 5'b11100: dout=32'b0001_0000_0000_0000_0000_0000_0000_0000;
	 5'b11101: dout=32'b0010_0000_0000_0000_0000_0000_0000_0000;
	 5'b11110: dout=32'b0100_0000_0000_0000_0000_0000_0000_0000;
	 5'b11111: dout=32'b1000_0000_0000_0000_0000_0000_0000_0000;
	endcase
  end
endmodule